module hi (
    a
);
    input a;
endmodule